module tof_top_test(


                    );
                    
endmodule